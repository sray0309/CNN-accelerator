

typedef enum {IDLE, LOAD, CONV, UPDATE} STATE;